library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library WORK;
use WORK.top_pack.all;


-------------------------------------------------------------------------------
package brick_position_pack is
-------------------------------------------------------------------------------

type t_init_pos_arr is array (0 to 3) of t_game_tile_pos;
type t_bricks_init_pos_arr is array (1 to C_NUM_OF_BRICKS) of t_init_pos_arr;
type t_next_pos_arr is array (0 to 3) of t_tile_pos;
type t_bricks_next_pos_arr is array (1 to C_NUM_OF_BRICKS) of t_next_pos_arr;

constant C_INIT_POS_ARR : t_bricks_init_pos_arr := (  
                               ( (5,1), (5,1), (5,0), (5,1) ), --Brick 1 (4 rotations)
                               ( (6,0), (5,2), (4,1), (5,0) ), --Brick 2
                               ( (5,0), (5,1), (5,0), (5,1) ), --Brick 3
                               ( (5,0), (5,1), (5,0), (5,1) ), --Brick 4
                               ( (5,0), (5,1), (5,0), (5,1) ), --Brick 5
                               ( (4,0), (5,0), (5,1), (5,2) ), --Brick 6
                               ( (6,0), (5,3), (6,0), (5,3) )  --Brick 7
                            );

constant C_NEXT_POS_ARR : t_bricks_next_pos_arr := (  
                                ( (35,16), (35,16), (35,15), (35,16) ), --Brick 1 (4 rotations)
                                ( (36,15), (35,17), (34,16), (35,15) ), --Brick 2
                                ( (35,15), (35,16), (35,15), (35,16) ), --Brick 3
                                ( (35,15), (35,16), (35,15), (35,16) ), --Brick 4
                                ( (35,15), (35,16), (35,15), (35,16) ), --Brick 5
                                ( (34,15), (35,15), (35,16), (35,17) ), --Brick 6
                                ( (36,15), (35,18), (36,15), (35,18) )  --Brick 7
                             );      

constant C_AI_NEXT_POS_ARR : t_bricks_next_pos_arr := (  
                                ( (41,10), (41,10), (41,9), (41,10) ), --Brick 1 (4 rotations)
                                ( (42,9), (41,11), (40,10), (41,9) ), --Brick 2
                                ( (41,9), (41,10), (41,9), (41,10) ), --Brick 3
                                ( (41,9), (41,10), (41,9), (41,10) ), --Brick 4
                                ( (41,9), (41,10), (41,9), (41,10) ), --Brick 5
                                ( (40,9), (41,9), (41,10), (41,11) ), --Brick 6
                                ( (42,9), (41,12), (42,9), (41,12) )  --Brick 7
                             ); 
--constant C_AI_NEXT_X_OFFSET : integer := 6;							 
--constant C_AI_NEXT_Y_OFFSET : integer := 4;							 
                             
type t_brick_move_pos is array (0 to 3) of t_pos_diff;                            
type t_brick_move_rec is record
    count           : integer range 1 to 4;
    elements_rw     : t_brick_move_pos;
    elements_del    : t_brick_move_pos;
end record;

type t_brick_move_map is array (0 to C_NUM_OF_MOVES-1) of t_brick_move_rec; -- moves
type t_brick_move_arr is array (0 to 3) of t_brick_move_map; -- 4 rot
type t_move_map is array (1 to C_NUM_OF_BRICKS) of t_brick_move_arr; -- 7 types 

constant C_MOVE_MAP : t_move_map :=
(
	(--1
		(
			(4,((0, 0), (-1, 0), (1, 0), (0, -1)),((0, 0), (-1, 0), (1, 0), (0, -1))),
			(3,((0, 1), (-1, 1), (1, 1), (0, 0)),((-1, 0), (1, 0), (0, -1), (0, 0))),
			(2,((-2, 0), (-1, -1), (0, 0), (0, 0)),((1, 0), (0, -1), (0, 0), (0, 0))),
			(2,((2, 0), (1, -1), (0, 0), (0, 0)),((-1, 0), (0, -1), (0, 0), (0, 0))),
			(1,((0, 1), (0, 0), (0, 0), (0, 0)),((-1, 0), (0, 0), (0, 0), (0, 0))),
			(1,((0, 1), (0, 0), (0, 0), (0, 0)),((1, 0), (0, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (1, 0), (0, -1), (0, 1)),((0, 0), (1, 0), (0, -1), (0, 1))),
			(2,((1, 1), (0, 2), (0, 0), (0, 0)),((1, 0), (0, -1), (0, 0), (0, 0))),
			(3,((-1, 0), (-1, -1), (-1, 1), (0, 0)),((1, 0), (0, -1), (0, 1), (0, 0))),
			(3,((2, 0), (1, -1), (1, 1), (0, 0)),((0, 0), (0, -1), (0, 1), (0, 0))),
			(1,((-1, 0), (0, 0), (0, 0), (0, 0)),((0, -1), (0, 0), (0, 0), (0, 0))),
			(1,((-1, 0), (0, 0), (0, 0), (0, 0)),((0, 1), (0, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (1, 0), (0, 1), (-1, 0)),((0, 0), (1, 0), (0, 1), (-1, 0))),
			(3,((1, 1), (0, 2), (-1, 1), (0, 0)),((0, 0), (1, 0), (-1, 0), (0, 0))),
			(2,((-1, 1), (-2, 0), (0, 0), (0, 0)),((1, 0), (0, 1), (0, 0), (0, 0))),
			(2,((2, 0), (1, 1), (0, 0), (0, 0)),((0, 1), (-1, 0), (0, 0), (0, 0))),
			(1,((0, -1), (0, 0), (0, 0), (0, 0)),((1, 0), (0, 0), (0, 0), (0, 0))),
			(1,((0, -1), (0, 0), (0, 0), (0, 0)),((-1, 0), (0, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, 1), (-1, 0), (0, -1)),((0, 0), (0, 1), (-1, 0), (0, -1))),
			(2,((0, 2), (-1, 1), (0, 0), (0, 0)),((-1, 0), (0, -1), (0, 0), (0, 0))),
			(3,((-1, 1), (-2, 0), (-1, -1), (0, 0)),((0, 0), (0, 1), (0, -1), (0, 0))),
			(3,((1, 0), (1, 1), (1, -1), (0, 0)),((0, 1), (-1, 0), (0, -1), (0, 0))),
			(1,((1, 0), (0, 0), (0, 0), (0, 0)),((0, 1), (0, 0), (0, 0), (0, 0))),
			(1,((1, 0), (0, 0), (0, 0), (0, 0)),((0, -1), (0, 0), (0, 0), (0, 0)))
		)
	),
	(--2
		(
			(4,((0, 0), (-1, 0), (-2, 0), (0, 1)),((0, 0), (-1, 0), (-2, 0), (0, 1))),
			(3,((-1, 1), (-2, 1), (0, 2), (0, 0)),((0, 0), (-1, 0), (-2, 0), (0, 0))),
			(2,((-3, 0), (-1, 1), (0, 0), (0, 0)),((0, 0), (0, 1), (0, 0), (0, 0))),
			(2,((1, 0), (1, 1), (0, 0), (0, 0)),((-2, 0), (0, 1), (0, 0), (0, 0))),
			(2,((0, -1), (0, -2), (0, 0), (0, 0)),((-2, 0), (0, 1), (0, 0), (0, 0))),
			(2,((0, 2), (1, 0), (0, 0), (0, 0)),((-1, 0), (-2, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (0, -2)),((0, 0), (-1, 0), (0, -1), (0, -2))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((-1, 0), (0, -2), (0, 0), (0, 0))),
			(3,((-2, 0), (-1, -1), (-1, -2), (0, 0)),((0, 0), (0, -1), (0, -2), (0, 0))),
			(3,((1, 0), (1, -1), (1, -2), (0, 0)),((-1, 0), (0, -1), (0, -2), (0, 0))),
			(2,((1, 0), (2, 0), (0, 0), (0, 0)),((-1, 0), (0, -2), (0, 0), (0, 0))),
			(2,((0, 1), (-2, 0), (0, 0), (0, 0)),((0, -1), (0, -2), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, -1), (1, 0), (2, 0)),((0, 0), (0, -1), (1, 0), (2, 0))),
			(3,((0, 1), (1, 1), (2, 1), (0, 0)),((0, -1), (1, 0), (2, 0), (0, 0))),
			(2,((-1, 0), (-1, -1), (0, 0), (0, 0)),((0, -1), (2, 0), (0, 0), (0, 0))),
			(2,((1, -1), (3, 0), (0, 0), (0, 0)),((0, 0), (0, -1), (0, 0), (0, 0))),
			(2,((0, 1), (0, 2), (0, 0), (0, 0)),((0, -1), (2, 0), (0, 0), (0, 0))),
			(2,((-1, 0), (0, -2), (0, 0), (0, 0)),((1, 0), (2, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (1, 0), (0, 1), (0, 2)),((0, 0), (1, 0), (0, 1), (0, 2))),
			(2,((1, 1), (0, 3), (0, 0), (0, 0)),((0, 0), (1, 0), (0, 0), (0, 0))),
			(3,((-1, 0), (-1, 1), (-1, 2), (0, 0)),((1, 0), (0, 1), (0, 2), (0, 0))),
			(3,((2, 0), (1, 1), (1, 2), (0, 0)),((0, 0), (0, 1), (0, 2), (0, 0))),
			(2,((-1, 0), (-2, 0), (0, 0), (0, 0)),((1, 0), (0, 2), (0, 0), (0, 0))),
			(2,((0, -1), (2, 0), (0, 0), (0, 0)),((0, 1), (0, 2), (0, 0), (0, 0)))
		)
	),
	(--3
		(
			(4,((0, 0), (-1, 0), (0, 1), (1, 1)),((0, 0), (-1, 0), (0, 1), (1, 1))),
			(3,((-1, 1), (0, 2), (1, 2), (0, 0)),((0, 0), (-1, 0), (1, 1), (0, 0))),
			(2,((-2, 0), (-1, 1), (0, 0), (0, 0)),((0, 0), (1, 1), (0, 0), (0, 0))),
			(2,((1, 0), (2, 1), (0, 0), (0, 0)),((-1, 0), (0, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, 1), (0, 0), (0, 0)),((0, 1), (1, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, 1), (0, 0), (0, 0)),((0, 1), (1, 1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (-1, 1)),((0, 0), (-1, 0), (0, -1), (-1, 1))),
			(2,((0, 1), (-1, 2), (0, 0), (0, 0)),((-1, 0), (0, -1), (0, 0), (0, 0))),
			(3,((-2, 0), (-1, -1), (-2, 1), (0, 0)),((0, 0), (0, -1), (-1, 1), (0, 0))),
			(3,((1, 0), (1, -1), (0, 1), (0, 0)),((-1, 0), (0, -1), (-1, 1), (0, 0))),
			(2,((0, 1), (1, 1), (0, 0), (0, 0)),((0, -1), (-1, 1), (0, 0), (0, 0))),
			(2,((0, 1), (1, 1), (0, 0), (0, 0)),((0, -1), (-1, 1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, 1), (1, 1)),((0, 0), (-1, 0), (0, 1), (1, 1))),
			(3,((-1, 1), (0, 2), (1, 2), (0, 0)),((0, 0), (-1, 0), (1, 1), (0, 0))),
			(2,((-2, 0), (-1, 1), (0, 0), (0, 0)),((0, 0), (1, 1), (0, 0), (0, 0))),
			(2,((1, 0), (2, 1), (0, 0), (0, 0)),((-1, 0), (0, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, 1), (0, 0), (0, 0)),((0, 1), (1, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, 1), (0, 0), (0, 0)),((0, 1), (1, 1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (-1, 1)),((0, 0), (-1, 0), (0, -1), (-1, 1))),
			(2,((0, 1), (-1, 2), (0, 0), (0, 0)),((-1, 0), (0, -1), (0, 0), (0, 0))),
			(3,((-2, 0), (-1, -1), (-2, 1), (0, 0)),((0, 0), (0, -1), (-1, 1), (0, 0))),
			(3,((1, 0), (1, -1), (0, 1), (0, 0)),((-1, 0), (0, -1), (-1, 1), (0, 0))),
			(2,((0, 1), (1, 1), (0, 0), (0, 0)),((0, -1), (-1, 1), (0, 0), (0, 0))),
			(2,((0, 1), (1, 1), (0, 0), (0, 0)),((0, -1), (-1, 1), (0, 0), (0, 0)))
		)
	),
	(--4
		(
			(4,((0, 0), (-1, 0), (-1, 1), (0, 1)),((0, 0), (-1, 0), (-1, 1), (0, 1))),
			(2,((-1, 2), (0, 2), (0, 0), (0, 0)),((0, 0), (-1, 0), (0, 0), (0, 0))),
			(2,((-2, 0), (-2, 1), (0, 0), (0, 0)),((0, 0), (0, 1), (0, 0), (0, 0))),
			(2,((1, 0), (1, 1), (0, 0), (0, 0)),((-1, 0), (-1, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, -1), (0, 0), (0, 0)),((-1, 1), (0, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, -1), (0, 0), (0, 0)),((-1, 1), (0, 1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (-1, -1)),((0, 0), (-1, 0), (0, -1), (-1, -1))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0))),
			(2,((-2, 0), (-2, -1), (0, 0), (0, 0)),((0, 0), (0, -1), (0, 0), (0, 0))),
			(2,((1, 0), (1, -1), (0, 0), (0, 0)),((-1, 0), (-1, -1), (0, 0), (0, 0))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (-1, 1), (0, 1)),((0, 0), (-1, 0), (-1, 1), (0, 1))),
			(2,((-1, 2), (0, 2), (0, 0), (0, 0)),((0, 0), (-1, 0), (0, 0), (0, 0))),
			(2,((-2, 0), (-2, 1), (0, 0), (0, 0)),((0, 0), (0, 1), (0, 0), (0, 0))),
			(2,((1, 0), (1, 1), (0, 0), (0, 0)),((-1, 0), (-1, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, -1), (0, 0), (0, 0)),((-1, 1), (0, 1), (0, 0), (0, 0))),
			(2,((0, -1), (-1, -1), (0, 0), (0, 0)),((-1, 1), (0, 1), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (-1, -1)),((0, 0), (-1, 0), (0, -1), (-1, -1))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0))),
			(2,((-2, 0), (-2, -1), (0, 0), (0, 0)),((0, 0), (0, -1), (0, 0), (0, 0))),
			(2,((1, 0), (1, -1), (0, 0), (0, 0)),((-1, 0), (-1, -1), (0, 0), (0, 0))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0))),
			(2,((0, 1), (-1, 1), (0, 0), (0, 0)),((0, -1), (-1, -1), (0, 0), (0, 0)))
		)
	),
	(--5
		(
			(4,((0, 0), (-1, 1), (0, 1), (1, 0)),((0, 0), (-1, 1), (0, 1), (1, 0))),
			(3,((-1, 2), (0, 2), (1, 1), (0, 0)),((0, 0), (-1, 1), (1, 0), (0, 0))),
			(2,((-1, 0), (-2, 1), (0, 0), (0, 0)),((0, 1), (1, 0), (0, 0), (0, 0))),
			(2,((1, 1), (2, 0), (0, 0), (0, 0)),((0, 0), (-1, 1), (0, 0), (0, 0))),
			(2,((-1, -1), (-1, 0), (0, 0), (0, 0)),((-1, 1), (1, 0), (0, 0), (0, 0))),
			(2,((-1, -1), (-1, 0), (0, 0), (0, 0)),((-1, 1), (1, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, 1), (-1, -1), (-1, 0)),((0, 0), (0, 1), (-1, -1), (-1, 0))),
			(2,((0, 2), (-1, 1), (0, 0), (0, 0)),((0, 0), (-1, -1), (0, 0), (0, 0))),
			(3,((-1, 1), (-2, -1), (-2, 0), (0, 0)),((0, 0), (0, 1), (-1, -1), (0, 0))),
			(3,((1, 0), (1, 1), (0, -1), (0, 0)),((0, 1), (-1, -1), (-1, 0), (0, 0))),
			(2,((1, 0), (-1, 1), (0, 0), (0, 0)),((-1, -1), (-1, 0), (0, 0), (0, 0))),
			(2,((1, 0), (-1, 1), (0, 0), (0, 0)),((-1, -1), (-1, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 1), (0, 1), (1, 0)),((0, 0), (-1, 1), (0, 1), (1, 0))),
			(3,((-1, 2), (0, 2), (1, 1), (0, 0)),((0, 0), (-1, 1), (1, 0), (0, 0))),
			(2,((-1, 0), (-2, 1), (0, 0), (0, 0)),((0, 1), (1, 0), (0, 0), (0, 0))),
			(2,((1, 1), (2, 0), (0, 0), (0, 0)),((0, 0), (-1, 1), (0, 0), (0, 0))),
			(2,((-1, -1), (-1, 0), (0, 0), (0, 0)),((-1, 1), (1, 0), (0, 0), (0, 0))),
			(2,((-1, -1), (-1, 0), (0, 0), (0, 0)),((-1, 1), (1, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, 1), (-1, -1), (-1, 0)),((0, 0), (0, 1), (-1, -1), (-1, 0))),
			(2,((0, 2), (-1, 1), (0, 0), (0, 0)),((0, 0), (-1, -1), (0, 0), (0, 0))),
			(3,((-1, 1), (-2, -1), (-2, 0), (0, 0)),((0, 0), (0, 1), (-1, -1), (0, 0))),
			(3,((1, 0), (1, 1), (0, -1), (0, 0)),((0, 1), (-1, -1), (-1, 0), (0, 0))),
			(2,((1, 0), (-1, 1), (0, 0), (0, 0)),((-1, -1), (-1, 0), (0, 0), (0, 0))),
			(2,((1, 0), (-1, 1), (0, 0), (0, 0)),((-1, -1), (-1, 0), (0, 0), (0, 0)))
		)
	),
	(--6
		(
			(4,((0, 0), (0, 1), (1, 0), (2, 0)),((0, 0), (0, 1), (1, 0), (2, 0))),
			(3,((0, 2), (1, 1), (2, 1), (0, 0)),((0, 0), (1, 0), (2, 0), (0, 0))),
			(2,((-1, 0), (-1, 1), (0, 0), (0, 0)),((0, 1), (2, 0), (0, 0), (0, 0))),
			(2,((1, 1), (3, 0), (0, 0), (0, 0)),((0, 0), (0, 1), (0, 0), (0, 0))),
			(2,((-1, 0), (0, 2), (0, 0), (0, 0)),((1, 0), (2, 0), (0, 0), (0, 0))),
			(2,((0, -1), (0, -2), (0, 0), (0, 0)),((0, 1), (2, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, 1), (-1, 0), (0, 2)),((0, 0), (0, 1), (-1, 0), (0, 2))),
			(2,((-1, 1), (0, 3), (0, 0), (0, 0)),((0, 0), (-1, 0), (0, 0), (0, 0))),
			(3,((-1, 1), (-2, 0), (-1, 2), (0, 0)),((0, 0), (0, 1), (0, 2), (0, 0))),
			(3,((1, 0), (1, 1), (1, 2), (0, 0)),((0, 1), (-1, 0), (0, 2), (0, 0))),
			(2,((0, -1), (-2, 0), (0, 0), (0, 0)),((0, 1), (0, 2), (0, 0), (0, 0))),
			(2,((1, 0), (2, 0), (0, 0), (0, 0)),((-1, 0), (0, 2), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (-1, 0), (0, -1), (-2, 0)),((0, 0), (-1, 0), (0, -1), (-2, 0))),
			(3,((0, 1), (-1, 1), (-2, 1), (0, 0)),((-1, 0), (0, -1), (-2, 0), (0, 0))),
			(2,((-1, -1), (-3, 0), (0, 0), (0, 0)),((0, 0), (0, -1), (0, 0), (0, 0))),
			(2,((1, 0), (1, -1), (0, 0), (0, 0)),((0, -1), (-2, 0), (0, 0), (0, 0))),
			(2,((1, 0), (0, -2), (0, 0), (0, 0)),((-1, 0), (-2, 0), (0, 0), (0, 0))),
			(2,((0, 1), (0, 2), (0, 0), (0, 0)),((0, -1), (-2, 0), (0, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, -1), (1, 0), (0, -2)),((0, 0), (0, -1), (1, 0), (0, -2))),
			(2,((0, 1), (1, 1), (0, 0), (0, 0)),((1, 0), (0, -2), (0, 0), (0, 0))),
			(3,((-1, 0), (-1, -1), (-1, -2), (0, 0)),((0, -1), (1, 0), (0, -2), (0, 0))),
			(3,((1, -1), (2, 0), (1, -2), (0, 0)),((0, 0), (0, -1), (0, -2), (0, 0))),
			(2,((0, 1), (2, 0), (0, 0), (0, 0)),((0, -1), (0, -2), (0, 0), (0, 0))),
			(2,((-1, 0), (-2, 0), (0, 0), (0, 0)),((1, 0), (0, -2), (0, 0), (0, 0)))
		)
	),
	(--7
		(
			(4,((0, 0), (-3, 0), (-2, 0), (-1, 0)),((0, 0), (-3, 0), (-2, 0), (-1, 0))),
			(4,((0, 1), (-3, 1), (-2, 1), (-1, 1)),((0, 0), (-3, 0), (-2, 0), (-1, 0))),
			(1,((-4, 0), (0, 0), (0, 0), (0, 0)),((0, 0), (0, 0), (0, 0), (0, 0))),
			(1,((1, 0), (0, 0), (0, 0), (0, 0)),((-3, 0), (0, 0), (0, 0), (0, 0))),
			(3,((0, -3), (0, -2), (0, -1), (0, 0)),((-3, 0), (-2, 0), (-1, 0), (0, 0))),
			(3,((0, -3), (0, -2), (0, -1), (0, 0)),((-3, 0), (-2, 0), (-1, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, -3), (0, -2), (0, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(1,((0, 1), (0, 0), (0, 0), (0, 0)),((0, -3), (0, 0), (0, 0), (0, 0))),
			(4,((-1, 0), (-1, -3), (-1, -2), (-1, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(4,((1, 0), (1, -3), (1, -2), (1, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(3,((-3, 0), (-2, 0), (-1, 0), (0, 0)),((0, -3), (0, -2), (0, -1), (0, 0))),
			(3,((-3, 0), (-2, 0), (-1, 0), (0, 0)),((0, -3), (0, -2), (0, -1), (0, 0)))
		),
		(
			(4,((0, 0), (-3, 0), (-2, 0), (-1, 0)),((0, 0), (-3, 0), (-2, 0), (-1, 0))),
			(4,((0, 1), (-3, 1), (-2, 1), (-1, 1)),((0, 0), (-3, 0), (-2, 0), (-1, 0))),
			(1,((-4, 0), (0, 0), (0, 0), (0, 0)),((0, 0), (0, 0), (0, 0), (0, 0))),
			(1,((1, 0), (0, 0), (0, 0), (0, 0)),((-3, 0), (0, 0), (0, 0), (0, 0))),
			(3,((0, -3), (0, -2), (0, -1), (0, 0)),((-3, 0), (-2, 0), (-1, 0), (0, 0))),
			(3,((0, -3), (0, -2), (0, -1), (0, 0)),((-3, 0), (-2, 0), (-1, 0), (0, 0)))
		),
		(
			(4,((0, 0), (0, -3), (0, -2), (0, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(1,((0, 1), (0, 0), (0, 0), (0, 0)),((0, -3), (0, 0), (0, 0), (0, 0))),
			(4,((-1, 0), (-1, -3), (-1, -2), (-1, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(4,((1, 0), (1, -3), (1, -2), (1, -1)),((0, 0), (0, -3), (0, -2), (0, -1))),
			(3,((-3, 0), (-2, 0), (-1, 0), (0, 0)),((0, -3), (0, -2), (0, -1), (0, 0))),
			(3,((-3, 0), (-2, 0), (-1, 0), (0, 0)),((0, -3), (0, -2), (0, -1), (0, 0)))
		)
	)
);





------------------------------------------------------------------------------- 
end brick_position_pack;
-------------------------------------------------------------------------------
